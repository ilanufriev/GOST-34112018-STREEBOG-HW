module strhw_p import strhw_common_types::*; #() (
    input  uint512            a_i,
    output uint512            result_o
  );

endmodule
