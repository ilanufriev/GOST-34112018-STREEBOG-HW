module tb #() ();

endmodule

