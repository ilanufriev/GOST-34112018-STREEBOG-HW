package strhw_common_types;

typedef enum logic[1:0] {
  CLEAR,
  BUSY,
  READY,
  DONE
} state_t;

typedef logic[511:0] uint512;
typedef logic[63:0]  uint64;
typedef logic[7:0]   uint8;
typedef logic[6:0]   uint7;

/* verilator lint_off UNUSEDPARAM */

// Huge constants (^ v ^ )
localparam uint512 INIT_VECTOR_512 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

localparam uint512 INIT_VECTOR_256 = 512'h01010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;

localparam C_SIZE = 12;

localparam BLOCK_SIZE = 64;

localparam ENABLE_DEBUG_OUTPUT = 1;

/* verilator lint_on UNUSEDPARAM */
endpackage
