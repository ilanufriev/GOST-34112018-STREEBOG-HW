package strhw_common_types;

typedef enum logic[1:0] {
  CLEAR,
  BUSY,
  READY,
  DONE
} state_t;

typedef logic[511:0] uint512;
typedef logic[5:0]   uint6;

// Huge constants (^ v ^ )

localparam uint512 INIT_VECTOR_512 = 512'h01010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;

localparam uint512 INIT_VECTOR_256 = 512'h01010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;

endpackage
