module tb #() ();

strhw_control_logic cl();

endmodule

