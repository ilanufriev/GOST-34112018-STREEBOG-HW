module strhw_sl import strhw_common_types::*; #() (
    input  uint512            a_i,
    output uint512            result_o
  );

endmodule
